`include "d_flip_flop_pulse_triggered.v"
