`include "half-adder.v"
