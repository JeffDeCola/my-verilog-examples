`include "decoder-3-8.v"
