`include "priority_arbiter.v"
