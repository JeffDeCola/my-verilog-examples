`include "jk_flip_flop_sync_clear.v"
