`include "single_port_ram_synchronous.v"
