`include "priority-arbiter.v"
