`include "mux-to-demux.v"

`include "../mux-4x1/mux-4x1.v"
`include "../demux-1x4/demux-1x4.v"