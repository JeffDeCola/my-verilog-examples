`include "jeff-74x151.v"
