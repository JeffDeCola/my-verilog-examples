`include "encoder-8-3.v"
