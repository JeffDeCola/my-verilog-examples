`include "xor2.v"
