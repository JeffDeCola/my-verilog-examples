`include "jeff_74x181.v"

`include "sections/input_section.v"
`include "sections/invert_m.v"
`include "sections/out_section_f3.v"
`include "sections/out_section_f2.v"
`include "sections/out_section_f1.v"
`include "sections/out_section_f0.v"
`include "sections/g_p_carry_section.v"
`include "sections/aeqb_section.v"
