`include "dual_port_ram_asynchronous.v"
