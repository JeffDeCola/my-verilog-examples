`include "encoder_8_3.v"
