`include "full_adder.v"
