`include "jeff_74x157.v"
