`include "simple_memory_using_1d_array.v"
