`include "jeff-74x161.v"

`include "sections/output-section.v"
`include "../../../basic-code/sequential-logic/jk-flip-flop/jk-flip-flop.v"