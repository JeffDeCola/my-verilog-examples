`timescale 1ns / 1ns
`include "jeff-74x181.v"

module jeff_74x181_tb;

// DATA TYPES - DECLAIR INPUTS AND OUTPUTS
reg  [3:0]  A, B, S;
reg         M, CI;
wire [3:0]  F;
wire        CO, AEQB, P, G;

// UUT
jeff_74x181 uut(
    .a3(A[3]), .a2(A[2]), .a1(A[1]), .a0(A[0]),
    .b3(B[3]), .b2(B[2]), .b1(B[1]), .b0(B[0]),
    .s3(S[3]), .s2(S[2]), .s1(S[1]), .s0(S[0]),
    .m(M), .ci(CI),
    .f3(F[3]), .f2(F[2]), .f1(F[1]), .f0(F[0]),
    .co(CO), .aeqb(AEQB), .p(P), .g(G)
);

// FILES
initial begin
    $dumpfile("jeff-74x181-tb.vcd");
    $dumpvars(0, jeff_74x181_tb);
end

// TESTCASE
initial begin
    $display("test start");
    S = 4'b0000; A = 4'b0000; B= 4'b0000;
    M = 0; CI = 0;

    // MODE = 1, CI = 0
    #15;  M = 1'b1; CI = 1'b0;
    #20;  S = 4'b0000; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0001; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0010; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0011; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0100; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0101; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0110; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0111; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1000; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1001; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1010; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1011; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1100; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1101; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1110; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1111; A = 4'b0000; B= 4'b0000; // F = ????
    
    // MODE = 0, CI = 0
    #20;  M = 1'b0; CI = 1'b0;
    #20;  S = 4'b0000; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0001; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0010; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0011; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0100; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0101; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0110; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0111; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1000; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1001; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1010; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1011; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1100; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1101; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1110; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1111; A = 4'b0000; B= 4'b0000; // F = ????

    // MODE = 0, CI = 1
    #20;  M = 1'b0; CI = 1'b1;
    #20;  S = 4'b0000; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0001; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0010; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0011; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0100; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0101; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0110; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b0111; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1000; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1001; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1010; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1011; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1100; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1101; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1110; A = 4'b0000; B= 4'b0000; // F = ????
    #20;  S = 4'b1111; A = 4'b0000; B= 4'b0000; // F = ????

    // DONE
    #20

    $display("test complete");
    $finish;
end

endmodule
