`include "jeff-74x157.v"
