`include "left_shift_register.v"
