`include "simple_8_bit_register.v"
