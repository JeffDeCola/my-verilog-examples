`include "simple-8-bit-register.v"
