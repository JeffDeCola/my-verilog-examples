`include "mux_to_demux.v"

`include "../mux_4x1/mux_4x1.v"
`include "../demux_1x4/demux_1x4.v"