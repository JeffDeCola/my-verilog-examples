`include "demux_1x4.v"
