`include "d-flip-flop.v"
