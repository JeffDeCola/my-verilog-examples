`include "t_flip_flop.v"
