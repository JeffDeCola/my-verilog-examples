// 4-input NAND gate
module and2(
    input           A, B,          //
    output          Y              //
);

// CONTINUOUS ASSIGNMENT STATEMENT
assign Y = A & B;

endmodule
