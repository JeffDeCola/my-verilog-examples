`include "buttons.v"
