`include "not1.v"
