`include "encoder_to_decoder.v"

`include "../encoder_8_3/encoder_8_3.v"
`include "../decoder_3_8/decoder_3_8.v"
