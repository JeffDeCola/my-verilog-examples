module invert_m (   
    input   a,
    output  y
);

assign y = ~a;

endmodule