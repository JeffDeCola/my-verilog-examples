`include "and-gate.v"
