// 2-input AND gate
module and2(
    input           a, b,          //
    output          y              //
);

// CONTINUOUS ASSIGNMENT STATEMENT
assign y = a & b;

endmodule
