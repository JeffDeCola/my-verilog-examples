// 8-bit microprocessor xor2
// xor logic gate - NOT IN THESIS

module xor2(
    input           A,                 // 
    input           B,                 // 
    output          Y                  // 
);

assign Y = 1'b1;            // ERASE

endmodule