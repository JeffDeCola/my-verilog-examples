`timescale 1ns / 100ps // time-unit = 1 ns, precision = 100 ps

// include files are in d_flip_flop_pos_edge_sync_en.vh

module D_FLIP_FLOP_POS_EDGE_SYNC_EN_TB ();

    // INPUT PROBES
    reg             EN;
    reg             D;

    // OUTPUT PROBES
    wire            Q_beh, QBAR_beh;

    // FOR TESTING  
    reg             CLK;
    reg [31:0]      VECTORCOUNT, ERRORS;
    reg             QEXPECTED;
    integer         FD, COUNT;
    reg [8*32-1:0]  COMMENT;

    // UNIT UNDER TEST (behavioral)
    d_flip_flop_pos_edge_sync_en_behavioral UUT_d_flip_flop_pos_edge_sync_en_behavioral(
        .clk(CLK),
        .en(EN),
        .d(D),
        .q(Q_beh), .qbar(QBAR_beh)
    );

    // SAVE EVERYTHING FROM TOP TB MODULE IN A DUMP FILE
    initial begin
        $dumpfile("d_flip_flop_pos_edge_sync_en_tb.vcd");
        $dumpvars(0, D_FLIP_FLOP_POS_EDGE_SYNC_EN_TB);
    end

    // CLK PERIOD
    localparam CLKPERIOD = 20;

    // CLK
    always begin
        #(CLKPERIOD/2) CLK = ~CLK;
    end

    // INITIALIZE TESTBENCH
    initial begin

        // OPEN VECTOR FILE - THROW AWAY FIRST LINE
        FD=$fopen("d_flip_flop_pos_edge_sync_en_tb.tv","r");
        COUNT = $fscanf(FD, "%s", COMMENT);
        // $display ("FIRST LINE IS: %s", COMMENT);

        // INIT TESTBENCH
        COUNT = $fscanf(FD, "%s %b %b %b", COMMENT, EN, D, QEXPECTED);
        CLK = 0;
        VECTORCOUNT = 1;
        ERRORS = 0;

        // DISPAY OUTPUT AND MONITOR
        $display();
        $display("TEST START --------------------------------");
        $display();
        $display("                               ");
        $display("                 | TIME(ns) | EN | D |  Q  |");
        $display("                 ---------------------------");
        // $monitor("%4d  %10s | %8d | %d  | %1d |  %1d  |", VECTORCOUNT, COMMENT, $time, EN, D, Q_beh);

    end

    // APPLY TEST VECTORS ON NEG EDGE CLK (ADD DELAY)
    always @(negedge CLK) begin

        // WAIT A BIT (AFTER CHECK)
        #5;

        // GET VECTORS FROM TB FILE
        COUNT = $fscanf(FD, "%s %b %b  %b", COMMENT, EN, D, QEXPECTED);

        // CHECK IF EOF - PRINT SUMMARY, CLOSE VECTOR FILE AND FINISH TB
        if (COUNT == -1) begin
            $fclose(FD);
            $display();
            $display(" VECTORS: %4d", VECTORCOUNT);
            $display("  ERRORS: %4d", ERRORS);
            $display();
            $display("TEST END ----------------------------------");
            $display();
            $finish;
        end

        // GET ANOTHER VECTOR
        VECTORCOUNT = VECTORCOUNT + 1;

    end

    // CHECK TEST VECTORS ON POS EGDE CLK
    always @(posedge CLK) begin

        // WAIT A BIT
        #5;

        // DISPLAY OUTPUT ON POS EDGE CLK
        $display("%4d  %10s | %8d | %d  | %1d |  %1d  |", VECTORCOUNT, COMMENT, $time, EN, D, Q_beh);

        // CHECK EACH VECTOR RESULT
        if (Q_beh !== QEXPECTED) begin
            $display("***ERROR (behavioral) - Expected Q = %b", QEXPECTED);
            ERRORS = ERRORS + 1;
        end

    end   

endmodule
