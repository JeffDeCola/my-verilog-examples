`include "demux-1x4.v"
