`include "simple_pipeline.v"
