`include "mealy_state_machine.v"
