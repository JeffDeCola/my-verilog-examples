`include "sr_latch.v"
