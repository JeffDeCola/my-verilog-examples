`include "decoder_3_8.v"
