`include "decoder_to_encoder.v"

`include "../decoder_3_8/decoder_3_8.v"
`include "../encoder_8_3/encoder_8_3.v"
