`include "sr_flip_flop.v"
