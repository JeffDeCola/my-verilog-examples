`include "dual_port_ram_synchronous.v"
