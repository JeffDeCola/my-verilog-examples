`include "nor2.v"
