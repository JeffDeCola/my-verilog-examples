module and_gate(
    x,
    y,
    xy
);

    input x, y;
    output xy;

    and(xy, x, y);

endmodule
