`include "pattern-recognition.v"
