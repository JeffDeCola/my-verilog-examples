// not1 gate
module not1 (
    input           a,             //
    output          y              //
);

// CONTINUOUS ASSIGNMENT STATEMENT
assign y = ~a;

endmodule
