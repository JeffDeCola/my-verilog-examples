`include "half_adder.v"
