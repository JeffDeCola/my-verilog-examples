// A synchronous fifo read pointer

module read_ptr (
    input             clk,              // Clock
    input             rst,              // Reset
    input             r_next,           // Read next
    output reg [3:0]  r_ptr);           // Read pointer

    // ALWAYS BLOCK with NON-BLOCKING PROCEDURAL ASSIGNMENT STATEMENT
    always @ (posedge clk) begin
        if (rst) begin
            r_ptr <= 3'b000;
        end else if (r_next) begin
            r_ptr <= r_ptr + 1;
        end else begin
            r_ptr <= r_ptr;
        end
    end

endmodule