`include "left-shift-register.v"
