`include "jk_flip_flop_pos_edge_sync_clear.v"
