`include "jk-flip-flop.v"
