`include "simple-memory-using-1d-array.v"
