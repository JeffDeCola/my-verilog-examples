`include "and_gates.v"
