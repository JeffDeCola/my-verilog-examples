`include "mux-4x1.v"
