`include "or2.v"
