`include "decoder-to-encoder.v"

`include "../decoder-3-8/decoder-3-8.v"
`include "../encoder-8-3/encoder-8-3.v"
