`include "mux_4x1.v"
