`include "jk_flip_flop.v"
