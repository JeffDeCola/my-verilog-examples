`include "fifo_synchronous.v"
