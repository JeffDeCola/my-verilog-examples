`include "and2.v"
