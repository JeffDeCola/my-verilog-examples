`include "moore_state_machine.v"
