`include "jeff_74x161.v"

`include "sections/output_section.v"
`include "../../../basic-code/sequential-logic//jk_flip_flop_pos_edge_sync_clear/jk_flip_flop_pos_edge_sync_clear.v"