module priority_arbitor(
    req_0,
    req_1,
    req_2,
    clk,
    rst,
    gnt_0,
    gnt_1,
    gnt_2,
);

    input req_0, req_1, req_2;
    input clk, rst;
    output gnt_0, gnt_1, gnt_2;

    wire req_0, req_1, req_2 ,clk;
    reg gnt_0, gnt_1, gnt_2;


endmodule
