`include "fifo_synchronous.v"
`include "../dual_port_ram_synchronous/dual_port_ram_synchronous.v"
