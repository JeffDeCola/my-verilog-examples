`include "d_flip_flop_pos_edge.v"
