// 2-input AND gate
module and2(
    input           A, B,          //
    output          Y              //
);

// CONTINUOUS ASSIGNMENT STATEMENT
assign y = a & b;

endmodule
