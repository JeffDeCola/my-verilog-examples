`include "d_flip_flop_pos_edge_sync_en.v"
