`include "full-adder.v"
