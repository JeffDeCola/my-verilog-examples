`include "d_flip_flop.v"
