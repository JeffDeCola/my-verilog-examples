`include "nand4.v"
