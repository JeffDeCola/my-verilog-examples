`include "simple-pipeline.v"
