`include "jeff-74x377.v"

`include "../../../basic-code/sequential-logic/d-flip-flop/d-flip-flop.v"
