`include "jeff_74x151.v"
